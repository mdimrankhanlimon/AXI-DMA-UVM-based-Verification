
interface clk_rst_interface;

    bit   CLK_1;
    bit   CLK_2;
    bit   clk;
    
    reg   RESET_1;
    reg   RESET_2;
    reg   rst_n;

endinterface   
