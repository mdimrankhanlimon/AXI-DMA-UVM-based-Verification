//`include "../../axi4_slave_uvc/axi4_slave_sequences/



