//`include "/home/cad_tech_02/LIMON/GITREPO/axi_dma_project/TB/clock_reset_uvc/clock_reset_sequences/sanity_simple_seq.sv"

`include "../../clock_reset_uvc/clock_reset_sequences/sanity_simple_seq.sv"


