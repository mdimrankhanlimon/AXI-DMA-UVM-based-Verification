
class clk_rst_agent_config extends uvm_object;
		`uvm_object_utils (clk_rst_agent_config)

		function new (string name = "clk_rst_agent_config");
				super.new(name);
		endfunction
endclass

