`define START_ADDR  32'h0000
`define END_ADDR    32'h2800
