////`include "base_test.sv"
`include "csr_wr_rd_test.sv"
`include "sanity_simple_test.sv"
`include "multiple_burst_transfer_test.sv"
`include "disable_descriptor_test.sv"
`include "error_response_test.sv"
`include "max_burst_configuration_test.sv"
`include "multiple_descriptor_configuration_test.sv"
`include "single_burst_transfer_test.sv"
`include "unaligned_source_transfer_test.sv"
`include "unaligned_destination_transfer_test.sv"
`include "abort_mid_transfer_test.sv"
`include "burst_exceeds_4k_boundary_test.sv"
`include "custom_test.sv"
`include "sample_sanity_test.sv"
`include "same_descriptor_multiple_configuration_test.sv"
